
module ROM(addr, data);
	input [31:0] addr;
	output reg [31:0] data;
	
	always @(*)
		case (addr[9:2])

			// Address:  0x00000000
// Instruct: 0x08000003		j Main
8'd0:  data = 32'b00001000000000000000000000000011;
8'd1:  data = 32'b00001000000000000000000000110101;
8'd2:  data = 32'b00001000000000000000000010101010;
8'd3:  data = 32'b00100000000011010000000000001000;
8'd4:  data = 32'b00100000000111010000001111111111;
8'd5:  data = 32'b00100000000010000000000001000000;
8'd6:  data = 32'b00111100000000100100000000000000;
8'd7:  data = 32'b00100000000010010000000000000011;
8'd8:  data = 32'b10101100010010010000000000100000;
8'd9:  data = 32'b10101100010000000000000000001000;
8'd10:  data = 32'b00100000000010010000001111101000;
8'd11:  data = 32'b00000000000010010100100000100010;
8'd12:  data = 32'b10101100010010010000000000000000;
8'd13:  data = 32'b00100000000010101111111111111111;
8'd14:  data = 32'b10101100010010100000000000000100;
8'd15:  data = 32'b00000001000000000000000000001000;
8'd16:  data = 32'b00100000000010100000000000000011;
8'd17:  data = 32'b10101100010010100000000000001000;
8'd18:  data = 32'b00000000000000001011000000100000;
8'd19:  data = 32'b00100000000100110000000000000010;
8'd20:  data = 32'b10001100010100000000000000100000;
8'd21:  data = 32'b00100000000101000000000000001000;
8'd22:  data = 32'b00000010100100001000100000100100;
8'd23:  data = 32'b00010110100100011111111111111100;
8'd24:  data = 32'b00010100000101100000000000000011;
8'd25:  data = 32'b10001100010001000000000000011100;
8'd26:  data = 32'b00100010110101100000000000000001;
8'd27:  data = 32'b00001000000000000000000000011110;
8'd28:  data = 32'b10001100010001010000000000011100;
8'd29:  data = 32'b00100010110101100000000000000001;
8'd30:  data = 32'b00000000000000001000100000100000;
8'd31:  data = 32'b00000010110100111000100000101010;
8'd32:  data = 32'b00010100000100011111111111110011;
8'd33:  data = 32'b00000000000000001011000000100000;
8'd34:  data = 32'b00001000000000000000000000100011;
8'd35:  data = 32'b00010100101001000000000000000010;
8'd36:  data = 32'b00000000100000001010100000100000;
8'd37:  data = 32'b00001000000000000000000000110001;
8'd38:  data = 32'b00000000100000001000100000100000;
8'd39:  data = 32'b00000000101000001001000000100000;
8'd40:  data = 32'b00000000000000001000000000100000;
8'd41:  data = 32'b00000010001100101000000000101010;
8'd42:  data = 32'b00010000000100000000000000000011;
8'd43:  data = 32'b00000010010000001010000000100000;
8'd44:  data = 32'b00000010001000001001000000100000;
8'd45:  data = 32'b00000010100000001000100000100000;
8'd46:  data = 32'b00000010001100101000100000100010;
8'd47:  data = 32'b00010110010100011111111111111000;
8'd48:  data = 32'b00000010001000001010100000100000;
8'd49:  data = 32'b10101100010101010000000000001100;
8'd50:  data = 32'b10101100010101010000000000011000;
8'd51:  data = 32'b00000010101000001010100000100000;
8'd52:  data = 32'b00001000000000000000000000010100;
8'd53:  data = 32'b00100000000010000000000000000001;
8'd54:  data = 32'b10101100010010000000000000001000;
8'd55:  data = 32'b00100000000010000000000000011000;
8'd56:  data = 32'b00000011101010001110100000100010;
8'd57:  data = 32'b10101111101100000000000000011000;
8'd58:  data = 32'b10101111101100010000000000010100;
8'd59:  data = 32'b10101111101100100000000000010000;
8'd60:  data = 32'b10101111101100110000000000001100;
8'd61:  data = 32'b10101111101101000000000000001000;
8'd62:  data = 32'b10101111101111110000000000000100;
8'd63:  data = 32'b00001100000000000000000001001110;
8'd64:  data = 32'b10001111101111110000000000000100;
8'd65:  data = 32'b10001111101101000000000000001000;
8'd66:  data = 32'b10001111101100110000000000001100;
8'd67:  data = 32'b10001111101100100000000000010000;
8'd68:  data = 32'b10001111101100010000000000010100;
8'd69:  data = 32'b10001111101100000000000000011000;
8'd70:  data = 32'b00100011101111010000000000011000;
8'd71:  data = 32'b10101100010000110000000000010100;
8'd72:  data = 32'b00100000000010010000000100110000;
8'd73:  data = 32'b00100000000010000000000000000011;
8'd74:  data = 32'b10101100010010000000000000001000;
8'd75:  data = 32'b00000000000000000100100000100000;
8'd76:  data = 32'b00100011010110101111111111111100;
8'd77:  data = 32'b00000011010000000000000000001000;
8'd78:  data = 32'b00000000000001000100011100000000;
8'd79:  data = 32'b00000000000010000100011100000010;
8'd80:  data = 32'b00000000000001000100100100000010;
8'd81:  data = 32'b00000000000001010101011100000000;
8'd82:  data = 32'b00000000000010100101011100000010;
8'd83:  data = 32'b00000000000001010101100100000010;
8'd84:  data = 32'b00100000000011100000000000001000;
8'd85:  data = 32'b00010001101011100000000000001001;
8'd86:  data = 32'b00000000000011100111000001000010;
8'd87:  data = 32'b00010001101011100000000000001011;
8'd88:  data = 32'b00000000000011100111000001000010;
8'd89:  data = 32'b00010001101011100000000000001101;
8'd90:  data = 32'b00000000000011100111000001000010;
8'd91:  data = 32'b00000000000011100001101000000000;
8'd92:  data = 32'b00000000000011010110100011000000;
8'd93:  data = 32'b00000000000010100111100000100000;
8'd94:  data = 32'b00001000000000000000000001101011;
8'd95:  data = 32'b00000000000011100001101000000000;
8'd96:  data = 32'b00000000000011010110100001000010;
8'd97:  data = 32'b00000000000010010111100000100000;
8'd98:  data = 32'b00001000000000000000000001101011;
8'd99:  data = 32'b00000000000011100001101000000000;
8'd100:  data = 32'b00000000000011010110100001000010;
8'd101:  data = 32'b00000000000010000111100000100000;
8'd102:  data = 32'b00001000000000000000000001101011;
8'd103:  data = 32'b00000000000011100001101000000000;
8'd104:  data = 32'b00000000000011010110100001000010;
8'd105:  data = 32'b00000000000010110111100000100000;
8'd106:  data = 32'b00001000000000000000000001101011;
8'd107:  data = 32'b00010000000011110000000000011110;
8'd108:  data = 32'b00100001111011111111111111111111;
8'd109:  data = 32'b00010000000011110000000000011110;
8'd110:  data = 32'b00100001111011111111111111111111;
8'd111:  data = 32'b00010000000011110000000000011110;
8'd112:  data = 32'b00100001111011111111111111111111;
8'd113:  data = 32'b00010000000011110000000000011110;
8'd114:  data = 32'b00100001111011111111111111111111;
8'd115:  data = 32'b00010000000011110000000000011110;
8'd116:  data = 32'b00100001111011111111111111111111;
8'd117:  data = 32'b00010000000011110000000000011110;
8'd118:  data = 32'b00100001111011111111111111111111;
8'd119:  data = 32'b00010000000011110000000000011110;
8'd120:  data = 32'b00100001111011111111111111111111;
8'd121:  data = 32'b00010000000011110000000000011110;
8'd122:  data = 32'b00100001111011111111111111111111;
8'd123:  data = 32'b00010000000011110000000000011110;
8'd124:  data = 32'b00100001111011111111111111111111;
8'd125:  data = 32'b00010000000011110000000000011110;
8'd126:  data = 32'b00100001111011111111111111111111;
8'd127:  data = 32'b00010000000011110000000000011110;
8'd128:  data = 32'b00100001111011111111111111111111;
8'd129:  data = 32'b00010000000011110000000000011110;
8'd130:  data = 32'b00100001111011111111111111111111;
8'd131:  data = 32'b00010000000011110000000000011110;
8'd132:  data = 32'b00100001111011111111111111111111;
8'd133:  data = 32'b00010000000011110000000000011110;
8'd134:  data = 32'b00100001111011111111111111111111;
8'd135:  data = 32'b00010000000011110000000000011110;
8'd136:  data = 32'b00100001111011111111111111111111;
8'd137:  data = 32'b00010000000011110000000000011110;
8'd138:  data = 32'b00100000011000110000000011000000;
8'd139:  data = 32'b00000011111000000000000000001000;
8'd140:  data = 32'b00100000011000110000000011111001;
8'd141:  data = 32'b00000011111000000000000000001000;
8'd142:  data = 32'b00100000011000110000000010100100;
8'd143:  data = 32'b00000011111000000000000000001000;
8'd144:  data = 32'b00100000011000110000000010110000;
8'd145:  data = 32'b00000011111000000000000000001000;
8'd146:  data = 32'b00100000011000110000000010011001;
8'd147:  data = 32'b00000011111000000000000000001000;
8'd148:  data = 32'b00100000011000110000000010010010;
8'd149:  data = 32'b00000011111000000000000000001000;
8'd150:  data = 32'b00100000011000110000000010000010;
8'd151:  data = 32'b00000011111000000000000000001000;
8'd152:  data = 32'b00100000011000110000000011111000;
8'd153:  data = 32'b00000011111000000000000000001000;
8'd154:  data = 32'b00100000011000110000000010000000;
8'd155:  data = 32'b00000011111000000000000000001000;
8'd156:  data = 32'b00100000011000110000000010010000;
8'd157:  data = 32'b00000011111000000000000000001000;
8'd158:  data = 32'b00100000011000110000000010001000;
8'd159:  data = 32'b00000011111000000000000000001000;
8'd160:  data = 32'b00100000011000110000000010000011;
8'd161:  data = 32'b00000011111000000000000000001000;
8'd162:  data = 32'b00100000011000110000000011000110;
8'd163:  data = 32'b00000011111000000000000000001000;
8'd164:  data = 32'b00100000011000110000000010100001;
8'd165:  data = 32'b00000011111000000000000000001000;
8'd166:  data = 32'b00100000011000110000000010000110;
8'd167:  data = 32'b00000011111000000000000000001000;
8'd168:  data = 32'b00100000011000110000000010001110;
8'd169:  data = 32'b00000011111000000000000000001000;
8'd170:  data = 32'b00000011010000000000000000001000;

			default: data = 32'h00000000;
		endcase
		
endmodule
